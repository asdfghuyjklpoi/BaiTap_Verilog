module A(input wire [2:0] X,output wire [2:0] Y);
assign Y = X - 3'b010;
endmodule