library verilog;
use verilog.vl_types.all;
entity tb_1 is
end tb_1;
